`timescale 1 ns / 100 ps

module CP4_processor_tb();

	reg clock, reset;
	wire [31:0] dmem_data_in, dmem_out;
	wire [11:0] dmem_address;

	CP4_processor_netid p(clock, reset, /*ps2_key_pressed, ps2_out, lcp.D_write, lcp.D_data,*/ dmem_data_in, dmem_address, dmem_out);

	initial
	begin
		clock = 0;
		reset = 0;
		
		@(negedge clock);
		
$monitor("<<<NEGEDGE>>>\nFETCH STAGE\ncurr_PC, %d, next_PC: %d\nchosen PC: %d, PC_jump: %b, PC_branch: %b, intialize PC: %b\np.F/D F instruction: %b\nDECODE STAGE\nopcode %b, rd %d, rs %d, rt %d, shamt %d, aluop %b, immediate %d, target %b\ninstrucion: add: %b, addi: %b, sub: %b, and: %b, or: %b, sll: %b, sra: %b, mul: %b, div: %b, sw: %b, lw: %b, j: %b, bne: %b, jal: %b, jr: %b, blt: %b, bex: %b, setx: %b\nreadAReg: %d, readBReg: %d, writeReg: %d\nEXECUTE STAGE\nDX_X_readA: %d, DX_X_readB: %d\nopcode %b, rd %d, rs %d, rt %d, shamt %d, real aluop: %b, aluop %b, immediate %d, target %b\ninstrucion: add: %d, addi: %d, sub: %d, and: %d, or: %d, sll: %d, sra: %d, mul: %d, div: %d, sw: %d, lw: %d, j: %d, bne: %d, jal: %d, jr: %d, blt: %d, bex: %d, setx: %d\n p.readAmemWrite: %d, p.readBmemWrite: %d, p.Amemequal: %d, p.Bmemequal: %d\np.readAwbWrite: %d, p.readBwbWrite: %d, p.Awbequal: %d, p.Bwbequal: %d\n\multdiv_status: %b, toggle_multdiv_status: %b, just_started: %b, multdiv_ready: %b, multdiv_ready,p.start_mul %b, p.start_div %b, p.my_multdiv.count %d\ndata_operandA: %d, data_operandB: %d\nX_alu_result: %d, X_multdiv_result: %d\not equal: %d, less than: %d\nMEMORY STAGE\nXM_M_op: %d, XM_M_readB: %d\nopcode %b, rd %d, rs %d, rt %d, shamt %d, aluop %b, immediate %d, target %b\ninstrucion: add: %d, addi: %d, sub: %d, and: %d, or: %d, sll: %d, sra: %d, mul: %d, div: %d, sw: %d, lw: %d, j: %d, bne: %d, jal: %d, jr: %d, blt: %d, bex: %d, setx: %d\ndmem_address %d, dmem_data_in: %d or %b, dmem_we: %d, dmem_out: %b, M_bex_taken: %b, curr rstatus: %d, next rstatus: %d\nWRITEBACK STAGE\nMW_W_op: %d, MW_W_data: %b\nopcode %b, rd %d, rs %d, rt %d, shamt %d, aluop %b, immediate %d, target %b\ninstrucion: add: %d, addi: %d, sub: %d, and: %d, or: %d, sll: %d, sra: %d, mul: %d, div: %d, sw: %d, lw: %d, j: %d, bne: %d, jal: %d, jr: %d, blt: %d, bex: %d, setx: %d\nreg_we: %b, write reg: %d, data %d\nregister[1]: %d\nregister[2]: %d\nregister[3]: %d\nregister[4]: %d\nregister[5]: %d\nregister[6]: %d\nregister[7]: %d\nregister[8]: %d\nregister[9]: %d\nregister[10]: %d\nregister[11]: %d\nregister[12]: %d\nregister[13]: %d\nregister[14]: %d\nregister[15]: %d\nregister[16]: %d\nregister[17]: %d\nregister[18]: %d\nregister[19]: %d\nregister[20]: %d\nregister[21]: %d\nregister[22]: %d\nregister[23]: %d\nregister[24]: %d\nregister[25]: %d\nregister[26]: %d\nregister[27]: %d\nregister[28]: %d\nregister[29]: %d\nregister[30]: %d\nregister[31]: %d\n p.PC_we %b,p.FD_we %b,p.DX_we %b,p.XM_we %b,p.MW_we %b",p.curr_PC, p.next_PC, p.imem_address, p.PC_jump, p.PC_branch, p.initialize_pc, p.FD_F_ir, p.D_op, p.D_rd, p.D_rs, p.D_rt, p.D_shamt, p.D_aluop, $signed(p.D_immediate), p.D_target, p.D_add,p.D_addi,p.D_sub,p.D_and,p.D_or, p.D_sll, p.D_sra, p.D_mul, p.D_div, p.D_sw, p.D_lw, p.D_j, p.D_bne, p.D_jal, p.D_jr, p.D_blt, p.D_bex, p.D_setx, p.regReadA, p.regReadB, p.regWrite, p.DX_X_readA,p.DX_X_readB,p.X_op, p.X_rd, p.X_rs, p.X_rt, p.X_shamt, p.alu_op, p.X_aluop, $signed(p.X_immediate), p.X_target, p.X_add,p.X_addi,p.X_sub,p.X_and,p.X_or, p.X_sll, p.X_sra, p.X_mul, p.X_div, p.X_sw, p.X_lw, p.X_j, p.X_bne, p.X_jal, p.X_jr, p.X_blt, p.X_bex, p.X_setx,p.readAmemWrite, p.readBmemWrite, p.Amemequal, p.Bmemequal,p.readAwbWrite, p.readBwbWrite, p.Awbequal, p.Bwbequal,p.multdiv_status, p.toggle_multdiv_status, p.just_started, p.multdiv_ready, p.start_mul, p.start_div, p.my_multdiv.count, $signed(p.data_operandA), $signed(p.data_operandB), p.X_alu_result, p.X_multdiv_result, p.X_isNotEqual, p.X_isLessThan, $signed(p.XM_M_op_result), $signed(p.XM_M_readB), p.M_op, p.M_rd, p.M_rs, p.M_rt, p.M_shamt, p.M_aluop, $signed(p.M_immediate), p.M_target, p.M_add,p.M_addi,p.M_sub,p.M_and,p.M_or, p.M_sll, p.M_sra, p.M_mul, p.M_div, p.M_sw, p.M_lw, p.M_j, p.M_bne, p.M_jal, p.M_jr, p.M_blt, p.M_bex, p.M_setx, p.dmem_address, $signed(p.dmem_data_in), p.dmem_data_in, p.dmem_we, p.MW_M_data_out, p.M_bex_taken, p.curr_rstatus_value, p.next_rstatus_value, $signed(p.MW_W_op_result),$signed(p.MW_W_data_out),p.W_op, p.W_rd, p.W_rs, p.W_rt, p.W_shamt, p.W_aluop, $signed(p.W_immediate), p.W_target, p.W_add,p.W_addi,p.W_sub,p.W_and,p.W_or, p.W_sll, p.W_sra, p.W_mul, p.W_div, p.W_sw, p.W_lw, p.W_j, p.W_bne, p.W_jal, p.W_jr, p.W_blt, p.W_bex, p.W_setx, p.reg_we,p.regWrite,$signed(p.regWrite_data),$signed(p.my_regfile.registeroutputdata[1]), $signed(p.my_regfile.registeroutputdata[2]), $signed(p.my_regfile.registeroutputdata[3]), $signed(p.my_regfile.registeroutputdata[4]), $signed(p.my_regfile.registeroutputdata[5]), $signed(p.my_regfile.registeroutputdata[6]), $signed(p.my_regfile.registeroutputdata[7]), $signed(p.my_regfile.registeroutputdata[8]), $signed(p.my_regfile.registeroutputdata[9]), $signed(p.my_regfile.registeroutputdata[10]), $signed(p.my_regfile.registeroutputdata[11]), $signed(p.my_regfile.registeroutputdata[12]), $signed(p.my_regfile.registeroutputdata[13]), $signed(p.my_regfile.registeroutputdata[14]), $signed(p.my_regfile.registeroutputdata[15]), $signed(p.my_regfile.registeroutputdata[16]), $signed(p.my_regfile.registeroutputdata[17]), $signed(p.my_regfile.registeroutputdata[18]), $signed(p.my_regfile.registeroutputdata[19]), $signed(p.my_regfile.registeroutputdata[20]), $signed(p.my_regfile.registeroutputdata[21]), $signed(p.my_regfile.registeroutputdata[22]), $signed(p.my_regfile.registeroutputdata[23]), $signed(p.my_regfile.registeroutputdata[24]), $signed(p.my_regfile.registeroutputdata[25]), $signed(p.my_regfile.registeroutputdata[26]), $signed(p.my_regfile.registeroutputdata[27]), $signed(p.my_regfile.registeroutputdata[28]), $signed(p.my_regfile.registeroutputdata[29]), $signed(p.my_regfile.registeroutputdata[30]), $signed(p.my_regfile.registeroutputdata[31]),p.PC_we,p.FD_we,p.DX_we,p.XM_we,p.MW_we);
	
		#2000
		$stop;

	end
	always
		#10 clock = ~clock;

endmodule