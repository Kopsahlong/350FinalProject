`timescale 1 ns / 100 ps

module processor_tb();

reg clock, reset, ps2_key_pressed, player1;
reg [7:0] ps2_out;

wire [31:0] dmem_data_in, dmem_out;

wire [11:0] dmem_address;
wire [9:0] score;


processor p(clock, reset, ps2_key_pressed, ps2_out, score, dmem_data_in, dmem_address, dmem_out, player1);



initial

begin
clock = 1'b1;
reset = 1'b0;
ps2_key_pressed = 1'b0;
player1 = 1'b1;
	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);

	

@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


@(posedge clock);
$display("<<<NEGEDGE>>>");
$display("p.PC_input, %d, p.PC_output: %d", p.PC_input, p.PC_output);
$display("p.instruction_FS: %b,\n p.opcode_FS: %b, p.ALU_op_FS %b, p.rd_FS: %d, p.rt_FS: %d, p.immediate_FS: %d, p.target_FS: %d", p.instruction_FS, p.opcode_FS, p.ALU_op_FS, p.rd_FS, p.rt_FS, p.immediate_FS, p.target_FS);
$display("p.instruction_DS: %b,\n p.opcode_DS: %b, p.ALU_op_DS %b, p.rd_DS: %d, p.rt_DS: %d, p.immediate_DS: %d, p.target_DS: %d", p.instruction_DS, p.opcode_DS, p.ALU_op_DS, p.rd_DS, p.rt_DS, p.immediate_DS, p.target_DS);
$display("p.instruction_XS: %b,\n p.opcode_XS: %b, p.ALU_op_XS %b, p.rd_XS: %d, p.rt_XS: %d, p.immediate_XS: %d, p.target_XS: %d", p.instruction_XS, p.opcode_XS, p.ALU_op_XS, p.rd_XS, p.rt_XS, p.immediate_XS, p.target_XS);
$display("p.instruction_MS: %b,\n p.opcode_MS: %b, p.ALU_op_MS %b, p.rd_MS: %d, p.rt_MS: %d, p.immediate_MS: %d, p.target_MS: %d", p.instruction_MS, p.opcode_MS, p.ALU_op_MS, p.rd_MS, p.rt_MS, p.immediate_MS, p.target_MS);
$display("p.instruction_WS: %b,\n p.opcode_WS: %b, p.ALU_op_WS %b, p.rd_WS: %d, p.rt_WS: %d, p.immediate_WS: %d, p.target_WS: %d", p.instruction_WS, p.opcode_WS, p.ALU_op_WS, p.rd_WS, p.rt_WS, p.immediate_WS, p.target_WS);
$display("score: %d", score);
$display("dmem_address: %b", p.dmem_address);
$display("dmem_data_in: %b", p.dmem_data_in);
$display("dmem_output_MS: %b", p.dmem_output_MS);
$display("p.regfile_WE: %b", p.regfile_WE);
$display("my_regfile.data_readReg_32b_1: %b", p.my_regfile.data_readReg_32b_1);
$display("my_regfile.data_readReg_32b_2: %b", p.my_regfile.data_readReg_32b_2);
$display("my_regfile.data_readReg_32b_3: %b", p.my_regfile.data_readReg_32b_3);
$display("my_regfile.data_readReg_32b_4: %b", p.my_regfile.data_readReg_32b_4);
$display("my_regfile.data_readReg_32b_5: %b", p.my_regfile.data_readReg_32b_5);
$display("my_regfile.data_readReg_32b_6: %b", p.my_regfile.data_readReg_32b_6);
$display("my_regfile.data_readReg_32b_7: %b", p.my_regfile.data_readReg_32b_7);
$display("my_regfile.data_readReg_32b_8: %b", p.my_regfile.data_readReg_32b_8);
$display("my_regfile.data_readReg_32b_9: %b", p.my_regfile.data_readReg_32b_9);
$display("my_regfile.data_readReg_32b_10: %b", p.my_regfile.data_readReg_32b_10);
$display("my_regfile.data_readReg_32b_11: %b", p.my_regfile.data_readReg_32b_11);
$display("my_regfile.data_readReg_32b_12: %b", p.my_regfile.data_readReg_32b_12);
$display("my_regfile.data_readReg_32b_13: %b", p.my_regfile.data_readReg_32b_13);
$display("my_regfile.data_readReg_32b_14: %b", p.my_regfile.data_readReg_32b_14);
$display("my_regfile.data_readReg_32b_15: %b", p.my_regfile.data_readReg_32b_15);
$display("my_regfile.data_readReg_32b_16: %b", p.my_regfile.data_readReg_32b_16);
$display("my_regfile.data_readReg_32b_17: %b", p.my_regfile.data_readReg_32b_17);
$display("my_regfile.data_readReg_32b_18: %b", p.my_regfile.data_readReg_32b_18);
$display("my_regfile.data_readReg_32b_19: %b", p.my_regfile.data_readReg_32b_19);
$display("my_regfile.data_readReg_32b_20: %b", p.my_regfile.data_readReg_32b_20);
$display("my_regfile.data_readReg_32b_21: %b", p.my_regfile.data_readReg_32b_21);
$display("my_regfile.data_readReg_32b_22: %b", p.my_regfile.data_readReg_32b_22);
$display("my_regfile.data_readReg_32b_23: %b", p.my_regfile.data_readReg_32b_23);
$display("my_regfile.data_readReg_32b_24: %b", p.my_regfile.data_readReg_32b_24);
$display("my_regfile.data_readReg_32b_25: %b", p.my_regfile.data_readReg_32b_25);
$display("my_regfile.data_readReg_32b_26: %b", p.my_regfile.data_readReg_32b_26);
$display("my_regfile.data_readReg_32b_27: %b", p.my_regfile.data_readReg_32b_27);
$display("my_regfile.data_readReg_32b_28: %b", p.my_regfile.data_readReg_32b_28);
$display("my_regfile.data_readReg_32b_29: %b", p.my_regfile.data_readReg_32b_29);
$display("my_regfile.data_readReg_32b_30: %b", p.my_regfile.data_readReg_32b_30);
$display("my_regfile.data_readReg_32b_31: %b", p.my_regfile.data_readReg_32b_31);


clock = 1'b0;

reset = 1'b0;

#300

$stop;

end



always

#10 clock = ~clock;

endmodule